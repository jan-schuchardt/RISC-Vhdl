----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:02:21 09/08/2016 
-- Design Name: 
-- Module Name:    BLOCKRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BLOCKRAM is
port(
		clk : in std_logic;
		rst : in std_logic;
		addr_in : in std_logic_vector(10 downto 0); --11 bit for adressing 8-bit cells
		data_in : in std_logic_vector(7 downto 0);
		data_out: out std_logic_vector(7 downto 0);
		write_enable : in std_logic
);

end BLOCKRAM;

architecture Behavioral of BLOCKRAM is

	type mem_t is array (0 to 2047) of std_logic_vector(7 downto 0);  -- 2048 cells with 8 bit
	signal cells : mem_t:=( --addi x1, x0, 0
"10010011","00000000","00000000","00000000",

--lui x1, 0x10000
"10110111","00000000","00000000","00010000",

--addi x2, x0, -1
"00010011","00000001","11110000","11111111",

--lui x3, 0x0F0F0
"10110111","00000001","00001111","00001111",

--addi x3, x3, 0x70F
"10010011","10000001","11110001","01110000",

--addi x3, x3, 0x700
"10010011","10000001","00000001","01110000",

--addi x3, x3, 0x100
"10010011","10000001","00000001","00010000",

--lui x4, 0xF0F0F
"00110111","11110010","11110000","11110000",

--addi x4, x4, 0xF0
"00010011","00000010","00000010","00001111",

--lui x5, 0x55555
"10110111","01010010","01010101","01010101",

--addi x5, x5, 0x555
"10010011","10000010","01010010","01010101",

--lui x6, 0x72AbE
"00110111","11100011","10101011","01110010",

--addi x6, x6, 0x9F0
"00010011","00000011","00000011","10011111",

--lui x7, 0xE7044
"10110111","01000011","00000100","11100111",

--addi x7, x7, 0xD71
"10010011","10000011","00010011","11010111",

--sw x1, x2, 0
"00100011","10100000","00100000","00000000",

--sw x1, x4, 8
"00100011","10100100","01000000","00000000",

--sw x1, x3, 4
"00100011","10100010","00110000","00000000",

--sw x1, x8, 12
"00100011","10100110","10000000","00000000",

--lw x10, x1, 8
"00000011","10100101","10000000","00000000",

--lw x8, x1, 0
"00000011","10100100","00000000","00000000",

--lw x11, x1, 12
"10000011","10100101","11000000","00000000",

--lw x9, x1, 4
"10000011","10100100","01000000","00000000",

--sw x1, x6, 0
"00100011","10100000","01100000","00000000",

--lw x15, x1, 12
"10000011","10100111","11000000","00000000",

--lw x13, x1, 4
"10000011","10100110","01000000","00000000",

--lw x12, x1, 0
"00000011","10100110","00000000","00000000",

--lw x14, x1, 8
"00000011","10100111","10000000","00000000",

--sw x1, x6, 5
"10100011","10100010","01100000","00000000",

--lw x16, x1, 0
"00000011","10101000","00000000","00000000",

--lw x19, x1, 12
"10000011","10101001","11000000","00000000",

--lw x17, x1, 4
"10000011","10101000","01000000","00000000",

--lw x18, x1, 8
"00000011","10101001","10000000","00000000",

--sh x1, x7, 8
"00100011","10010100","01110000","00000000",

--lw x21, x1, 5
"10000011","10101010","01010000","00000000",

--lw x20, x1, 1
"00000011","10101010","00010000","00000000",

--lw x23, x1, 13
"10000011","10101011","11010000","00000000",

--lw x22, x1, 9
"00000011","10101011","10010000","00000000",

--sh x1, x7, 11
"10100011","10010101","01110000","00000000",

--lw x26, x1, 10
"00000011","10101101","10100000","00000000",

--lw x27, x1, 14
"10000011","10101101","11100000","00000000",

--lb x24, x1, 2
"00000011","10001100","00100000","00000000",

--lh x25, x1, 6
"10000011","10011100","01100000","00000000",

--sb x1, x7, 14
"00100011","10000111","01110000","00000000",

--lb x28, x1, 3
"00000011","10001110","00110000","00000000",

--lw x31, x1, 15
"10000011","10101111","11110000","00000000",

--lh x29, x1, 7
"10000011","10011110","01110000","00000000",

--lw x30, x1, 11
"00000011","10101111","10110000","00000000",

others=>(others=>'0')

	);
	
	attribute ram_style: string;
	attribute ram_style of cells : signal is "block";
	
begin
	

	process(clk) begin
	
		
		
		if rising_edge(clk) then
		
			if rst = '0' then
			--No reset -> standard dual-port usage
				if write_enable = '1'then
					cells(to_integer(unsigned(addr_in))) <= data_in;
				end if;
				data_out <= cells(to_integer(unsigned(addr_in)));
			
			end if;
			
			
			
			
		end if;
			
	end process;

end Behavioral;
