----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    11:02:21 09/08/2016 
-- Design Name: 
-- Module Name:    BLOCKRAM - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity BLOCKRAM is
port(
		clk : in std_logic;
		rst : in std_logic;
		addr_in : in std_logic_vector(10 downto 0); --11 bit for adressing 8-bit cells
		data_in : in std_logic_vector(7 downto 0);
		data_out: out std_logic_vector(7 downto 0);
		write_enable : in std_logic
);

end BLOCKRAM;

architecture Behavioral of BLOCKRAM is

	type mem_t is array (0 to 2047) of std_logic_vector(7 downto 0);  -- 2048 cells with 8 bit
	signal cells : mem_t:= (--addi x2, x2, 0x400
"00010011","00000001","00000001","01000000",

--addi x2, x2, 0x400
"00010011","00000001","00000001","01000000",

--jal x0, main
"01101111","00000000","01000000","00101100",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x2D2D2D2D
"00101101","00101101","00101101","00101101",

--dw 0x00007C7C
"01111100","01111100","00000000","00000000",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x7C7C0000
"00000000","00000000","01111100","01111100",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x00007C7C
"01111100","01111100","00000000","00000000",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x7C7C0000
"00000000","00000000","01111100","01111100",

--dw 0x0000005C
"01011100","00000000","00000000","00000000",

--dw 0x2F2F2F00
"00000000","00101111","00101111","00101111",

--dw 0x2F5C0000
"00000000","00000000","01011100","00101111",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x5C2F0000
"00000000","00000000","00101111","01011100",

--dw 0x00000000
"00000000","00000000","00000000","00000000",

--dw 0x0000002F
"00101111","00000000","00000000","00000000",

--dw 0x00005C00
"00000000","01011100","00000000","00000000",

--dw 0x2D2D2800
"00000000","00101000","00101101","00101101",

--dw 0x00000029
"00101001","00000000","00000000","00000000",

--dw 0x00000028
"00101000","00000000","00000000","00000000",

--dw 0x00002900
"00000000","00101001","00000000","00000000",

--dw 0x00000028
"00101000","00000000","00000000","00000000",

--dw 0x00002900
"00000000","00101001","00000000","00000000",

--dw 0x2D2D2800
"00000000","00101000","00101101","00101101",

--dw 0x00000029
"00101001","00000000","00000000","00000000",

--dw 0x65697053
"01010011","01110000","01101001","01100101",

--dw 0x2072656C
"01101100","01100101","01110010","00100000",

--dw 0x73692031
"00110001","00100000","01101001","01110011",

--dw 0x6D612074
"01110100","00100000","01100001","01101101",

--dw 0x67755A20
"00100000","01011010","01110101","01100111",

--dw 0x0000002E
"00101110","00000000","00000000","00000000",

--dw 0x65697053
"01010011","01110000","01101001","01100101",

--dw 0x2072656C
"01101100","01100101","01110010","00100000",

--dw 0x65672031
"00110001","00100000","01100111","01100101",

--dw 0x6E6E6977
"01110111","01101001","01101110","01101110",

--dw 0x00002E74
"01110100","00101110","00000000","00000000",

--addi x2, x2, -8
"00010011","00000001","10000001","11111111",

--sw x2, x1, 0
"00100011","00100000","00010001","00000000",

--sw x2, x3, 4
"00100011","00100010","00110001","00000000",

--addi x3, x0, 15
"10010011","00000001","11110000","00000000",

--blt x3, x0, end_setup_border
"01100011","11000100","00000001","00000100",

--addi x18, x0, vborder
"00010011","00001001","11000000","00000010",

--slli x27, x3, 6
"10010011","10011101","01100001","00000000",

--lui x19, 0x20000
"10110111","00001001","00000000","00100000",

--addi x19, x19, 64
"10010011","10001001","00001001","00000100",

--add x19, x19, x27
"10110011","10001001","10111001","00000001",

--addi x26, x0, 15
"00010011","00001101","11110000","00000000",

--beq x3, x26, phbord
"01100011","10001100","10100001","00000001",

--addi x26, x0, 10
"00010011","00001101","10100000","00000000",

--beq x3, x26, phbord
"01100011","10001000","10100001","00000001",

--addi x26, x0, 5
"00010011","00001101","01010000","00000000",

--beq x3, x26, phbord
"01100011","10000100","10100001","00000001",

--bne x3, x0, wboard
"01100011","10010100","00000001","00000000",

--addi x18, x0, hborder
"00010011","00001001","11000000","00000000",

--addi x20, x0, 32
"00010011","00001010","00000000","00000010",

--jal x1, memcpy
"11101111","00000000","01000000","00110110",

--addi x3, x3, -1
"10010011","10000001","11110001","11111111",

--jal x0, setup_border_loop
"01101111","11110000","11011111","11111011",

--lw x1, x2, 0
"10000011","00100000","00000001","00000000",

--lw x3, x2, 4
"10000011","00100001","01000001","00000000",

--addi x2, x2, 8
"00010011","00000001","10000001","00000000",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--addi x2, x2, -16
"00010011","00000001","00000001","11111111",

--sw x2, x1, 0
"00100011","00100000","00010001","00000000",

--sw x2, x3, 4
"00100011","00100010","00110001","00000000",

--sw x2, x4, 8
"00100011","00100100","01000001","00000000",

--sw x2, x5, 12
"00100011","00100110","01010001","00000000",

--addi x26, x0, 10
"00010011","00001101","10100000","00000000",

--mul x26, x26, x18
"00110011","00001101","00101101","00000011",

--addi x26, x26, 3
"00010011","00001101","00111101","00000000",

--addi x27, x0, 5
"10010011","00001101","01010000","00000000",

--mul x19, x19, x27
"10110011","10001001","10111001","00000011",

--addi x19, x19, 1
"10010011","10001001","00011001","00000000",

--slli x19, x19, 6
"10010011","10011001","01101001","00000000",

--add x3, x19, x26
"10110011","10000001","10101001","00000001",

--addi x5, x0, 4
"10010011","00000010","01000000","00000000",

--addi x4, x0, cross
"00010011","00000010","11000000","00000100",

--beq x20, x0, do_print_element
"01100011","00000100","00001010","00000000",

--addi x4, x0, dot
"00010011","00000010","11000000","00000110",

--beq x5, x0, end_print_element
"01100011","10000110","00000010","00000010",

--addi x18, x4, 0
"00010011","00001001","00000010","00000000",

--lui x19, 0x20000
"10110111","00001001","00000000","00100000",

--addi x19, x19, 64
"10010011","10001001","00001001","00000100",

--add x19, x19, x3
"10110011","10001001","00111001","00000000",

--addi x20, x0, 6
"00010011","00001010","01100000","00000000",

--jal x1, memcpy
"11101111","00000000","11000000","00101110",

--addi x5, x5, -1
"10010011","10000010","11110010","11111111",

--addi x4, x4, 8
"00010011","00000010","10000010","00000000",

--addi x3, x3, 64
"10010011","10000001","00000001","00000100",

--jal x0, do_print_element
"01101111","11110000","10011111","11111101",

--lw x1, x2, 0
"10000011","00100000","00000001","00000000",

--lw x3, x2, 4
"10000011","00100001","01000001","00000000",

--lw x4, x2, 8
"00000011","00100010","10000001","00000000",

--lw x5, x2, 12
"10000011","00100010","11000001","00000000",

--addi x2, x2, 16
"00010011","00000001","00000001","00000001",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--addi x26, x0, 10
"00010011","00001101","10100000","00000000",

--mul x26, x26, x18
"00110011","00001101","00101101","00000011",

--addi x27, x0, 5
"10010011","00001101","01010000","00000000",

--mul x27, x27, x19
"10110011","10001101","00111101","00000011",

--addi x27, x27, 1
"10010011","10001101","00011101","00000000",

--slli x27, x27, 6
"10010011","10011101","01101101","00000000",

--lui x28, 0x20000
"00110111","00001110","00000000","00100000",

--addi x28, x28, 64
"00010011","00001110","00001110","00000100",

--add x26, x26, x27
"00110011","00001101","10111101","00000001",

--add x26, x26, x28
"00110011","00001101","11001101","00000001",

--addi x29, x0, 4
"10010011","00001110","01000000","00000000",

--addi x28, x0, 0x0
"00010011","00001110","00000000","00000000",

--beq x20, x0, do_cursor_set_active
"01100011","00000100","00001010","00000000",

--addi x28, x0, 0x2A
"00010011","00001110","10100000","00000010",

--beq x29, x0, end_cursor_set_active
"01100011","10001100","00001110","00000000",

--sb x26, x28, 2
"00100011","00000001","11001101","00000001",

--sb x26, x28, 9
"10100011","00000100","11001101","00000001",

--addi x26, x26, 64
"00010011","00001101","00001101","00000100",

--addi x29, x29, -1
"10010011","10001110","11111110","11111111",

--jal x0, do_cursor_set_active
"01101111","11110000","11011111","11111110",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x26, 0x30000
"00110111","00001101","00000000","00110000",

--lh x27, x26, 0
"10000011","00011101","00001101","00000000",

--srli x27, x27, 7
"10010011","11011101","01111101","00000000",

--andi x27, x27, 0x1F
"10010011","11111101","11111101","00000001",

--lh x28, x26, 0
"00000011","00011110","00001101","00000000",

--srli x28, x28, 7
"00010011","01011110","01111110","00000000",

--andi x28, x28, 0x1F
"00010011","01111110","11111110","00000001",

--addi x30, x28, 0
"00010011","00001111","00001110","00000000",

--xor x28, x28, x27
"00110011","01001110","10111110","00000001",

--and x28, x28, x27
"00110011","01111110","10111110","00000001",

--addi x27, x30, 0
"10010011","00001101","00001111","00000000",

--beq x28, x0, key_release_wait
"11100011","00000010","00001110","11111110",

--addi x18, x0, 0
"00010011","00001001","00000000","00000000",

--addi x29, x0, 1
"10010011","00001110","00010000","00000000",

--beq x28, x29, end_key_release
"01100011","00001000","11011110","00000001",

--srli x28, x28, 1
"00010011","01011110","00011110","00000000",

--addi x18, x18, 1
"00010011","00001001","00011001","00000000",

--jal x0, key_release_shift_result
"01101111","11110000","01011111","11111111",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x26, 0x10000
"00110111","00001101","00000000","00010000",

--sb x26, x18, 0
"00100011","00000000","00101101","00000001",

--lui x26, 0x30000
"00110111","00001101","00000000","00110000",

--lui x28, 0x20000
"00110111","00001110","00000000","00100000",

--addi x28, x28, 0x440
"00010011","00001110","00001110","01000100",

--addi x27, x0, 0
"10010011","00001101","00000000","00000000",

--addi x29, x0, 0x31
"10010011","00001110","00010000","00000011",

--beq x18, x0, set_turn_set_led
"01100011","00000110","00001001","00000000",

--addi x27, x0, 1
"10010011","00001101","00010000","00000000",

--addi x29, x29, 1
"10010011","10001110","00011110","00000000",

--sb x26, x27, 2
"00100011","00000001","10111101","00000001",

--sb x28, x29, 8
"00100011","00000100","11011110","00000001",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x26, 0x10000
"00110111","00001101","00000000","00010000",

--lb x18, x26, 0
"00000011","00001001","00001101","00000000",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x26, 0x10000
"00110111","00001101","00000000","00010000",

--addi x27, x0, -4
"10010011","00001101","11000000","11111111",

--sw x26, x27, 4
"00100011","00100010","10111101","00000001",

--sw x26, x27, 8
"00100011","00100100","10111101","00000001",

--sb x26, x27, 12
"00100011","00000110","10111101","00000001",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x26, 0x10000
"00110111","00001101","00000000","00010000",

--addi x27, x0, 3
"10010011","00001101","00110000","00000000",

--mul x27, x19, x27
"10110011","10001101","10111001","00000011",

--add x27, x27, x18
"10110011","10001101","00101101","00000001",

--add x27, x27, x26
"10110011","10001101","10101101","00000001",

--lb x26, x27, 4
"00000011","10001101","01001101","00000000",

--addi x18, x0, 0
"00010011","00001001","00000000","00000000",

--bge x26, x0, end_matrix_can_place
"01100011","01010110","00001101","00000000",

--sb x27, x20, 4
"00100011","10000010","01001101","00000001",

--addi x18, x0, 1
"00010011","00001001","00010000","00000000",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--lui x3, 0x20000
"10110111","00000001","00000000","00100000",

--addi x3, x3, 0x440
"10010011","10000001","00000001","01000100",

--addi x18, x0, 0
"00010011","00001001","00000000","00000000",

--addi x19, x3, 0
"10010011","10001001","00000001","00000000",

--addi x20, x0, 64
"00010011","00001010","00000000","00000100",

--jal x1, memfill
"11101111","00000000","10000000","00011010",

--addi x19, x3, 0
"10010011","10001001","00000001","00000000",

--addi x18, x0, str_player_turn
"00010011","00001001","11000000","00001000",

--addi x20, x0, 24
"00010011","00001010","10000000","00000001",

--jal x1, memcpy
"11101111","00000000","10000000","00010111",

--addi x18, x0, 0
"00010011","00001001","00000000","00000000",

--jal x1, set_turn
"11101111","11110000","00011111","11110101",

--jal x1, matrix_init
"11101111","11110000","11011111","11111000",

--addi x3, x0, 1
"10010011","00000001","00010000","00000000",

--addi x4, x0, 1
"00010011","00000010","00010000","00000000",

--jal x1, setup_border
"11101111","11110000","00011111","11011011",

--addi x18, x3, 0
"00010011","10001001","00000001","00000000",

--addi x19, x4, 0
"10010011","00001001","00000010","00000000",

--addi x20, x0, 1
"00010011","00001010","00010000","00000000",

--jal x1, cursor_set_active
"11101111","11110000","00011111","11101001",

--jal x1, key_release
"11101111","11110000","00011111","11101110",

--addi x26, x0, 4
"00010011","00001101","01000000","00000000",

--addi x6, x18, 0
"00010011","00000011","00001001","00000000",

--beq x6, x26, request_place_element
"01100011","00001100","10100011","00000011",

--addi x18, x3, 0
"00010011","10001001","00000001","00000000",

--addi x19, x4, 0
"10010011","00001001","00000010","00000000",

--addi x20, x0, 0
"00010011","00001010","00000000","00000000",

--jal x1, cursor_set_active
"11101111","11110000","00011111","11100111",

--addi x27, x0, 3
"10010011","00001101","00110000","00000000",

--addi x26, x0, 1
"00010011","00001101","00010000","00000000",

--beq x6, x26, btn_north
"01100011","00001110","10100011","00000111",

--addi x26, x0, 2
"00010011","00001101","00100000","00000000",

--beq x6, x26, btn_south
"01100011","00000000","10100011","00001001",

--addi x26, x0, 3
"00010011","00001101","00110000","00000000",

--beq x6, x26, btn_west
"01100011","00001000","10100011","00001001",

--beq x6, x0, btn_east
"01100011","00000000","00000011","00001000",

--jal x0, idle_loop
"01101111","11110000","00011111","11111100",

--jal x1, get_turn
"11101111","11110000","11011111","11110001",

--addi x5, x18, 0
"10010011","00000010","00001001","00000000",

--addi x18, x3, 0
"00010011","10001001","00000001","00000000",

--addi x19, x4, 0
"10010011","00001001","00000010","00000000",

--addi x20, x5, 0
"00010011","10001010","00000010","00000000",

--jal x1, matrix_place_if_possible
"11101111","11110000","11011111","11110010",

--beq x18, x0, idle_loop
"11100011","00000010","00001001","11111010",

--addi x18, x3, 0
"00010011","10001001","00000001","00000000",

--addi x19, x4, 0
"10010011","00001001","00000010","00000000",

--addi x20, x5, 0
"00010011","10001010","00000010","00000000",

--jal x1, print_element
"11101111","11110000","10011111","11011001",

--xori x18, x5, 1
"00010011","11001001","00010010","00000000",

--jal x1, set_turn
"11101111","11110000","10011111","11101011",

--jal x0, idle_loop
"01101111","11110000","10011111","11111000",

--blt x18, x0, idle_loop
"11100011","01000010","00001001","11111000",

--addi x3, x18, 0
"10010011","00000001","00001001","00000000",

--addi x18, x0, str_player_won
"00010011","00001001","01000000","00001010",

--lui x19, 0x20000
"10110111","00001001","00000000","00100000",

--addi x19, x19, 0x440
"10010011","10001001","00001001","01000100",

--addi x20, x0, 20
"00010011","00001010","01000000","00000001",

--jal x1, memcpy
"11101111","00000000","10000000","00001011",

--lui x19 0x20000
"10110111","00001001","00000000","00100000",

--addi x19, x19, 0x440
"10010011","10001001","00001001","01000100",

--sb x19, x3, 8
"00100011","10000100","00111001","00000000",

--addi x4, x4, 2
"00010011","00000010","00100010","00000000",

--rem x4, x4, x27
"00110011","01100010","10110010","00000011",

--jal x0, cursor_update
"01101111","00000000","01000000","00000010",

--addi x4, x4, 1
"00010011","00000010","00010010","00000000",

--rem x4, x4, x27
"00110011","01100010","10110010","00000011",

--jal x0, cursor_update
"01101111","00000000","10000000","00000001",

--addi x3, x3, 1
"10010011","10000001","00010001","00000000",

--rem x3, x3, x27
"10110011","11100001","10110001","00000011",

--jal x0, cursor_update
"01101111","00000000","11000000","00000000",

--addi x3, x3, 2
"10010011","10000001","00100001","00000000",

--rem x3, x3, x27
"10110011","11100001","10110001","00000011",

--addi x18, x3, 0
"00010011","10001001","00000001","00000000",

--addi x19, x4, 0
"10010011","00001001","00000010","00000000",

--addi x20, x0, 1
"00010011","00001010","00010000","00000000",

--jal x1, cursor_set_active
"11101111","11110000","00011111","11011011",

--jal x0, idle_loop
"01101111","11110000","00011111","11110010",

--lui x26, 0x10000
"00110111","00001101","00000000","00010000",

--addi x27, x26, 0
"10010011","00001101","00001101","00000000",

--addi x28, x0, 2
"00010011","00001110","00100000","00000000",

--addi x18, x0, -1
"00010011","00001001","11110000","11111111",

--blt x28, x0, end_player_won_hv_loop
"01100011","01001010","00001110","00000100",

--addi x29, x0, 3
"10010011","00001110","00110000","00000000",

--addi x30, x0, 0
"00010011","00001111","00000000","00000000",

--addi x31, x0, 0
"10010011","00001111","00000000","00000000",

--add x19, x26, x28
"10110011","00001001","11001101","00000001",

--addi x20, x0, 3
"00010011","00001010","00110000","00000000",

--mul x20, x28, x20
"00110011","00001010","01001110","00000011",

--add x20, x26, x20
"00110011","00001010","01001101","00000001",

--beq x29, x0, end_player_won_inner
"01100011","10001110","00001110","00000000",

--lb x21, x19, 4
"10000011","10001010","01001001","00000000",

--add x31, x31, x21
"10110011","10001111","01011111","00000001",

--lb x21, x20, 4
"10000011","00001010","01001010","00000000",

--add x30, x30, x21
"00110011","00001111","01011111","00000001",

--addi x20, x20, -1
"00010011","00001010","11111010","11111111",

--jal x0, player_won_inner
"01101111","11110000","10011111","11111110",

--addi x28, x28, -1
"00010011","00001110","11111110","11111111",

--bge x30, x0, player_won_hsum
"01100011","01010110","00001111","00000000",

--blt x31, x0, player_won_hv_loop
"11100011","11001110","00001111","11111010",

--addi x30, x31, 0
"00010011","10001111","00001111","00000000",

--addi x19, x0, 3
"10010011","00001001","00110000","00000000",

--div x18, x30, x19
"00110011","01001001","00111111","00000011",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--beq x20, x0, end_memcpy
"01100011","00001110","00001010","00000000",

--lb x26, x18, 0
"00000011","00001101","00001001","00000000",

--sb x19, x26, 0
"00100011","10000000","10101001","00000001",

--addi x18, x18, 1
"00010011","00001001","00011001","00000000",

--addi x19, x19, 1
"10010011","10001001","00011001","00000000",

--addi x20, x20, -1
"00010011","00001010","11111010","11111111",

--jal x0, memcpy
"01101111","11110000","10011111","11111110",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

--beq x20, x0, end_memfill
"01100011","00001010","00001010","00000000",

--sb x19, x18, 0
"00100011","10000000","00101001","00000001",

--addi x19, x19, 1
"10010011","10001001","00011001","00000000",

--addi x20, x20, -1
"00010011","00001010","11111010","11111111",

--jal x0, memfill
"01101111","11110000","00011111","11111111",

--jalr x0, x1, 0
"01100111","10000000","00000000","00000000",

others=>(others=>'0')




	);
	
	attribute ram_style: string;
	attribute ram_style of cells : signal is "block";
	
begin
	

	process(clk) begin
	
		
		
		if rising_edge(clk) then
		
			if rst = '0' then
			--No reset -> standard dual-port usage
				if write_enable = '1'then
					cells(to_integer(unsigned(addr_in))) <= data_in;
				end if;
				data_out <= cells(to_integer(unsigned(addr_in)));
			
			end if;
			
			
			
			
		end if;
			
	end process;

end Behavioral;
