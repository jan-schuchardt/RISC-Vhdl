-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: Franz
-- 
-- Create Date:    10/11/2016 22:40:10
-- Project Name:   Ascii
-- Module Name:    Ascii.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity Ascii is
--   port( );
end Ascii;

architecture arq1 of Ascii is
begin

end arq1;
